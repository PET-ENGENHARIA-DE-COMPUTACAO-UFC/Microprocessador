module shift_left8b(input[7:0]a, output[7:0]y);
assign y = a << 1'b1;
endmodule